module main

fn main() {
	mut a := 5
	a = 3
	println(a)
}
