module main

fn main() {
	a := fn (n u32) u32 {
		return n + 1
	}

	println(a(3))
}
