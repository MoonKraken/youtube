module main

import src.some_module

fn main() {
	println(a.add(1, 3))
}
