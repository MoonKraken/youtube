module main

fn main() {
	mut a := 2 + 2
	a = 5
	println(a)
}
