module main

fn some_fun(n int) int {
	return n + 1
}

fn main() {
	println(some_fun(2))
}
